//-------------------------------------------------------------------------
//                                                                       --
//                                                                       --
//      For use with ECE 385 Lab 62                                       --
//      UIUC ECE Department                                              --
//-------------------------------------------------------------------------


module lab62 (

      ///////// Clocks /////////
      input     MAX10_CLK1_50, 

      ///////// KEY /////////
      input    [ 1: 0]   KEY,

      ///////// SW /////////
      input    [ 9: 0]   SW,

      ///////// LEDR /////////
      output   [ 9: 0]   LEDR,

      ///////// HEX /////////
      output   [ 7: 0]   HEX0,
      output   [ 7: 0]   HEX1,
      output   [ 7: 0]   HEX2,
      output   [ 7: 0]   HEX3,
      output   [ 7: 0]   HEX4,
      output   [ 7: 0]   HEX5,

      ///////// SDRAM /////////
      output             DRAM_CLK,
      output             DRAM_CKE,
      output   [12: 0]   DRAM_ADDR,
      output   [ 1: 0]   DRAM_BA,
      inout    [15: 0]   DRAM_DQ,
      output             DRAM_LDQM,
      output             DRAM_UDQM,
      output             DRAM_CS_N,
      output             DRAM_WE_N,
      output             DRAM_CAS_N,
      output             DRAM_RAS_N,

      ///////// VGA /////////
      output             VGA_HS,
      output             VGA_VS,
      output   [ 7: 0]   VGA_R,
      output   [ 7: 0]   VGA_G,
      output   [ 7: 0]   VGA_B,


      ///////// ARDUINO /////////
      inout    [15: 0]   ARDUINO_IO,
      inout              ARDUINO_RESET_N 

);




logic Run_h, Reset_h, vssig, blank, sync, VGA_Clk;


//=======================================================
//  REG/WIRE declarations
//=======================================================
	logic SPI0_CS_N, SPI0_SCLK, SPI0_MISO, SPI0_MOSI, USB_GPX, USB_IRQ, USB_RST;
	logic [3:0] hex_num_4, hex_num_3, hex_num_1, hex_num_0; //4 bit input hex digits
	logic [1:0] signs;
	logic [1:0] hundreds;
	logic [9:0] drawxsig, drawysig, ballxsig, ballysig, ballsizesig;
	logic [7:0] red, blue, green;
	logic [7:0] keycode;

//=======================================================
//  Structural coding
//=======================================================
	assign ARDUINO_IO[10] = SPI0_CS_N;
	assign ARDUINO_IO[13] = SPI0_SCLK;
	assign ARDUINO_IO[11] = SPI0_MOSI;
	assign ARDUINO_IO[12] = 1'bZ;
	assign SPI0_MISO = ARDUINO_IO[12];
	
	assign ARDUINO_IO[9] = 1'bZ; 
	assign USB_IRQ = ARDUINO_IO[9];
		
	//Assignments specific to Circuits At Home UHS_20
	assign ARDUINO_RESET_N = USB_RST;
	assign ARDUINO_IO[7] = USB_RST;//USB reset 
	assign ARDUINO_IO[8] = 1'bZ; //this is GPX (set to input)
	assign USB_GPX = 1'b0;//GPX is not needed for standard USB host - set to 0 to prevent interrupt
	
	//Assign uSD CS to '1' to prevent uSD card from interfering with USB Host (if uSD card is plugged in)
	assign ARDUINO_IO[6] = 1'b1;
	
	//HEX drivers to convert numbers to HEX output
	HexDriver hex_driver4 (hex_num_4, HEX4[6:0]);
	assign HEX4[7] = 1'b1;
	
	HexDriver hex_driver3 (hex_num_3, HEX3[6:0]);
	assign HEX3[7] = 1'b1;
	
	HexDriver hex_driver1 (hex_num_1, HEX1[6:0]);
	assign HEX1[7] = 1'b1;
	
	HexDriver hex_driver0 (hex_num_0, HEX0[6:0]);
	assign HEX0[7] = 1'b1;
	
	//fill in the hundreds digit as well as the negative sign
	assign HEX5 = {1'b1, ~signs[1], 3'b111, ~hundreds[1], ~hundreds[1], 1'b1};
	assign HEX2 = {1'b1, ~signs[0], 3'b111, ~hundreds[0], ~hundreds[0], 1'b1};
	
	
	//Assign one button to reset
	assign {Reset_h}=~ (KEY[0]);
	
	//Assign another button to run
	assign {Run_h}=~ (KEY[1]);

	//Our A/D converter is only 12 bit
	assign VGA_R = red[7:4];
	assign VGA_B = blue[7:4];
	assign VGA_G = green[7:4];
	
	
	lab62_soc u0 (
		.clk_clk                           (MAX10_CLK1_50),  //clk.clk
		.reset_reset_n                     (1'b1),           //reset.reset_n
		.altpll_0_locked_conduit_export    (),               //altpll_0_locked_conduit.export
		.altpll_0_phasedone_conduit_export (),               //altpll_0_phasedone_conduit.export
		.altpll_0_areset_conduit_export    (),               //altpll_0_areset_conduit.export
		.key_external_connection_export    (KEY),            //key_external_connection.export

		//SDRAM
		.sdram_clk_clk(DRAM_CLK),                            //clk_sdram.clk
		.sdram_wire_addr(DRAM_ADDR),                         //sdram_wire.addr
		.sdram_wire_ba(DRAM_BA),                             //.ba
		.sdram_wire_cas_n(DRAM_CAS_N),                       //.cas_n
		.sdram_wire_cke(DRAM_CKE),                           //.cke
		.sdram_wire_cs_n(DRAM_CS_N),                         //.cs_n
		.sdram_wire_dq(DRAM_DQ),                             //.dq
		.sdram_wire_dqm({DRAM_UDQM,DRAM_LDQM}),              //.dqm
		.sdram_wire_ras_n(DRAM_RAS_N),                       //.ras_n
		.sdram_wire_we_n(DRAM_WE_N),                         //.we_n

		//USB SPI	
		.spi0_SS_n(SPI0_CS_N),
		.spi0_MOSI(SPI0_MOSI),
		.spi0_MISO(SPI0_MISO),
		.spi0_SCLK(SPI0_SCLK),
		
		//USB GPIO
		.usb_rst_export(USB_RST),
		.usb_irq_export(USB_IRQ),
		.usb_gpx_export(USB_GPX),
		
		//LEDs and HEX
		.hex_digits_export({hex_num_4, hex_num_3, hex_num_1, hex_num_0}),
		.leds_export({hundreds, signs, LEDR}),
		.keycode_export(keycode)
		
	 );

//other necesssary REG/WIRE
	logic game_over, game_reset, touching, shape_reset, stopxleft, stopxright;
	logic [1:0] screen_state, rotation;
	logic [2:0] shape_num, next_shape, next_shape2, key_state;
	logic [9:0] shape_size_x, shape_size_y, shape_x, shape_y;
	logic [19:0][9:0][3:0] PMO;
	logic [13:0] Score;
	logic [4:0] thousand_digit, hundred_digit, ten_digit, single_digit;
	
	/*
	assign shape_num = 3'd2;
	assign next_shape = 3'd2;
	assign next_shape2 = 3'd2;
	*/
	
//module instatiation
	vga_controller VGA(.Clk(MAX10_CLK1_50), .Reset(Reset_h), .hs(VGA_HS), .vs(VGA_VS),
							 .pixel_clk(VGA_Clk), .blank(blank), .sync(sync),
							 .DrawX(drawxsig), .DrawY(drawysig) );
	
//wait state for pressing a key on keyboard
	keywait keys(.Clk(MAX10_CLK1_50), .Reset(Reset_h), 
					 .keycode(keycode), 
					 .key(key_state));	

//FSM for handling rotation of a piece
	rotating rotate(.Clk(MAX10_CLK1_50), .Reset(Reset_h), 
						 .keycode(keycode), 
						 .rotation(rotation));

//FSM for determining what the screen is meant to be displaying
	screen gameplay(.Clk(MAX10_CLK1_50), .Reset(Reset_h), 
						 .game_over(game_over), 
						 .keycode(keycode),
						 .game_reset(game_reset), 
						 .screen_state(screen_state));

//bag of 7 random generator
	random_piece RNG(.Clk(MAX10_CLK1_50), .Reset(Reset_h), 
						  .shape_reset(shape_reset), .touching(touching), 
						  .shape_num(shape_num), .next_shape(next_shape), .next_shape2(next_shape2),
						  .game_over(game_over));

//dimension determination of a piece in a given rotation
	block_shape shape_n_rot(.shape_num(shape_num), .rotation(rotation), 
									.shape_size_x(shape_size_x), .shape_size_y(shape_size_y));
	
//datapath to control what is goin on
	datapath Tetris(.Clk(MAX10_CLK1_50), .Reset(Reset_h), .game_reset(game_reset), .frame_clk(VGA_VS),
						 .shape_num(shape_num), .rotation(rotation),  .keypress(key_state), .state(screen_state), 
						 .shape_size_x(shape_size_x), .shape_size_y(shape_size_y), .shape_x(shape_x), .shape_y(shape_y), 
						 .PixelMapOut(PMO), .shape_reset(shape_reset), .touching(touching), .theScore(Score),
						 .game_over(game_over), .stopxleft(stopxleft), .stopxright(stopxright));

//displaying the current acticity to the screen
	color_mapper color(.DrawX(drawxsig), .DrawY(drawysig), 
							 .shape_size_x(shape_size_x), .shape_size_y(shape_size_y), .shape_x(shape_x), .shape_y(shape_y), 
							 .keycode(keycode), 
							 .shape_num(shape_num), .next_shape(next_shape), .next_shape2(next_shape2), 
							 .game_state(screen_state), .rotation(rotation), .PixelMapOut(PMO),
							 .thousand(thousand_digit), .hundred(hundred_digit), .ten(ten_digit), .ones(single_digit),
							 .Red(red), .Green(green), .Blue(blue));
							 
	Score_Board game_score (.Reset(Reset_h),
									.Score(Score),
									.thousands(thousand_digit),
									.hundreds(hundred_digit),
									.tens(ten_digit),
									.ones(single_digit));
	

//	ball blocks(.Reset(Reset_h), .frame_clk(VGA_VS), .keycode(keycode), .Run(Run_h),
//					.BallX(ballxsig), .BallY(ballysig), .BallS(ballsizesig) );
endmodule
