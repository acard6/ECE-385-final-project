//each block is 4x4 chunck where each chuck is 4 bits wide
//each bit represetns a single pixel on the screen

module sprites_table_block( output logic [3:0][3:0][3:0] I_block_UB,
									 output logic [3:0][3:0][3:0] O_block_UB,
									 output logic [3:0][3:0][3:0] J_block_UB,
									 output logic [3:0][3:0][3:0] T_block_UB,
									 output logic [3:0][3:0][3:0] L_block_UB,
									 output logic [3:0][3:0][3:0] S_block_UB,
									 output logic [3:0][3:0][3:0] Z_block_UB);
	always_comb	
	 begin
	 //this maps the blocks of a tetromino to their respective color
		I_block_UB = '{
		'{1,1,1,1},
		'{1,1,1,1},
		'{1,1,1,1},
		'{1,1,1,1}
		};
		
		O_block_UB = '{
		'{2,2,2,2},
		'{2,2,2,2},
		'{2,2,2,2},
		'{2,2,2,2}
		};
		
		J_block_UB = '{
		'{3,3,3,3},
		'{3,3,3,3},
		'{3,3,3,3},
		'{3,3,3,3}
		};
		
		L_block_UB = ' {
		'{4,4,4,4},
		'{4,4,4,4},
		'{4,4,4,4},
		'{4,4,4,4}
		};

		S_block_UB = '{
		'{5,5,5,5},
		'{5,5,5,5},
		'{5,5,5,5},
		'{5,5,5,5}
		};
		
		Z_block_UB = '{
		'{6,6,6,6},
		'{6,6,6,6},
		'{6,6,6,6},
		'{6,6,6,6}
		};
		
		T_block_UB = '{
		'{7,7,7,7},
		'{7,7,7,7},
		'{7,7,7,7},
		'{7,7,7,7}
		};
	 end	
endmodule 

module sprite_table_font(
					 output logic [10:0][24:0][3:0]	game_over,
					 output logic [4:0][39:0][3:0] 	TETRIS_h,
					 output logic [3:0][15:0][3:0] 	I_block_h,
					 output logic [15:0][3:0][3:0] 	I_block_v,
					 output logic [7:0][7:0][3:0] 	O_block,
					 output logic [7:0][11:0][3:0]	J_block_0,
					 output logic [11:0][7:0][3:0]	J_block_1,
					 output logic [7:0][11:0][3:0]	J_block_2,
					 output logic [11:0][7:0][3:0] 	J_block_3,
					 output logic [7:0][11:0][3:0] 	T_block_0,
					 output logic [11:0][7:0][3:0] 	T_block_1,
					 output logic [7:0][11:0][3:0] 	T_block_2,
					 output logic [11:0][7:0][3:0] 	T_block_3,
					 output logic [7:0][11:0][3:0] 	L_block_0,
					 output logic [11:0][7:0][3:0] 	L_block_1,
					 output logic [7:0][11:0][3:0] 	L_block_2,
					 output logic [11:0][7:0][3:0] 	L_block_3,
					 output logic [7:0][11:0][3:0] 	S_block_0,
					 output logic [11:0][7:0][3:0] 	S_block_1,
					 output logic [7:0][11:0][3:0] 	Z_block_0,
					 output logic [11:0][7:0][3:0] 	Z_block_1,
					 output logic [4:0][28:0][3:0] SCORE_Letters,
					 output logic [4:0][4:0][3:0] zero,
					 output logic [4:0][4:0][3:0] one,
					 output logic [4:0][4:0][3:0] two,
					 output logic [4:0][4:0][3:0] three,
					 output logic [4:0][4:0][3:0] four,
					 output logic [4:0][4:0][3:0] five,
					 output logic [4:0][4:0][3:0] six,
					 output logic [4:0][4:0][3:0] seven,
					 output logic [4:0][4:0][3:0] eight,
					 output logic [4:0][4:0][3:0] nine);
	
	always_comb
	 begin
		
		I_block_h = '{
		'{1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1},
		'{1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1},
		'{1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1},
		'{1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1}};
		
		I_block_v = '{
		'{1,1,1,1},
		'{1,1,1,1},
		'{1,1,1,1},
		'{1,1,1,1},
		'{1,1,1,1},
		'{1,1,1,1},
		'{1,1,1,1},
		'{1,1,1,1},
		'{1,1,1,1},
		'{1,1,1,1},
		'{1,1,1,1},
		'{1,1,1,1},
		'{1,1,1,1},
		'{1,1,1,1},
		'{1,1,1,1},
		'{1,1,1,1}};


		O_block = '{
		'{2,2,2,2,2,2,2,2},
		'{2,2,2,2,2,2,2,2},
		'{2,2,2,2,2,2,2,2},
		'{2,2,2,2,2,2,2,2},
		'{2,2,2,2,2,2,2,2},
		'{2,2,2,2,2,2,2,2},
		'{2,2,2,2,2,2,2,2},
		'{2,2,2,2,2,2,2,2}};
		
		J_block_0 = '{
		'{3,3,3,3,3,3,3,3,3,3,3,3},
		'{3,3,3,3,3,3,3,3,3,3,3,3},
		'{3,3,3,3,3,3,3,3,3,3,3,3},
		'{3,3,3,3,3,3,3,3,3,3,3,3},
		'{0,0,0,0,0,0,0,0,3,3,3,3},
		'{0,0,0,0,0,0,0,0,3,3,3,3},
		'{0,0,0,0,0,0,0,0,3,3,3,3},
		'{0,0,0,0,0,0,0,0,3,3,3,3}};
		
		J_block_1 = '{
		'{0,0,0,0,3,3,3,3},
		'{0,0,0,0,3,3,3,3},
		'{0,0,0,0,3,3,3,3},
		'{0,0,0,0,3,3,3,3},
		'{0,0,0,0,3,3,3,3},
		'{0,0,0,0,3,3,3,3},
		'{0,0,0,0,3,3,3,3},
		'{0,0,0,0,3,3,3,3},
		'{3,3,3,3,3,3,3,3},
		'{3,3,3,3,3,3,3,3},
		'{3,3,3,3,3,3,3,3},
		'{3,3,3,3,3,3,3,3}};
		
		J_block_2 = '{
		'{3,3,3,3,0,0,0,0,0,0,0,0},
		'{3,3,3,3,0,0,0,0,0,0,0,0},
		'{3,3,3,3,0,0,0,0,0,0,0,0},
		'{3,3,3,3,0,0,0,0,0,0,0,0},
		'{3,3,3,3,3,3,3,3,3,3,3,3},
		'{3,3,3,3,3,3,3,3,3,3,3,3},
		'{3,3,3,3,3,3,3,3,3,3,3,3},
		'{3,3,3,3,3,3,3,3,3,3,3,3}};
		
		J_block_3 = '{
		'{3,3,3,3,3,3,3,3},
		'{3,3,3,3,3,3,3,3},
		'{3,3,3,3,3,3,3,3},
		'{3,3,3,3,3,3,3,3},
		'{3,3,3,3,0,0,0,0},
		'{3,3,3,3,0,0,0,0},
		'{3,3,3,3,0,0,0,0},
		'{3,3,3,3,0,0,0,0},
		'{3,3,3,3,0,0,0,0},
		'{3,3,3,3,0,0,0,0},
		'{3,3,3,3,0,0,0,0},
		'{3,3,3,3,0,0,0,0}};
		
		L_block_0 = ' {
		'{4,4,4,4,4,4,4,4,4,4,4,4},
		'{4,4,4,4,4,4,4,4,4,4,4,4},
		'{4,4,4,4,4,4,4,4,4,4,4,4},
		'{4,4,4,4,4,4,4,4,4,4,4,4},
		'{4,4,4,4,0,0,0,0,0,0,0,0},
		'{4,4,4,4,0,0,0,0,0,0,0,0},
		'{4,4,4,4,0,0,0,0,0,0,0,0},
		'{4,4,4,4,0,0,0,0,0,0,0,0}};
		
		L_block_1 = ' {
		'{4,4,4,4,4,4,4,4},
		'{4,4,4,4,4,4,4,4},
		'{4,4,4,4,4,4,4,4},
		'{4,4,4,4,4,4,4,4},
		'{0,0,0,0,4,4,4,4},
		'{0,0,0,0,4,4,4,4},
		'{0,0,0,0,4,4,4,4},
		'{0,0,0,0,4,4,4,4},
		'{0,0,0,0,4,4,4,4},
		'{0,0,0,0,4,4,4,4},
		'{0,0,0,0,4,4,4,4},
		'{0,0,0,0,4,4,4,4}};
		
		L_block_2 = ' {
		'{0,0,0,0,0,0,0,0,4,4,4,4},
		'{0,0,0,0,0,0,0,0,4,4,4,4},
		'{0,0,0,0,0,0,0,0,4,4,4,4},
		'{0,0,0,0,0,0,0,0,4,4,4,4},
		'{4,4,4,4,4,4,4,4,4,4,4,4},
		'{4,4,4,4,4,4,4,4,4,4,4,4},
		'{4,4,4,4,4,4,4,4,4,4,4,4},
		'{4,4,4,4,4,4,4,4,4,4,4,4}};
		
		L_block_3 = ' {
		'{4,4,4,4,0,0,0,0},
		'{4,4,4,4,0,0,0,0},
		'{4,4,4,4,0,0,0,0},
		'{4,4,4,4,0,0,0,0},
		'{4,4,4,4,0,0,0,0},
		'{4,4,4,4,0,0,0,0},
		'{4,4,4,4,0,0,0,0},
		'{4,4,4,4,0,0,0,0},
		'{4,4,4,4,4,4,4,4},
		'{4,4,4,4,4,4,4,4},
		'{4,4,4,4,4,4,4,4},
		'{4,4,4,4,4,4,4,4}};
		
		S_block_0 = '{
		'{0,0,0,0,6,6,6,6,6,6,6,6},
		'{0,0,0,0,6,6,6,6,6,6,6,6},
		'{0,0,0,0,6,6,6,6,6,6,6,6},
		'{0,0,0,0,6,6,6,6,6,6,6,6},
		'{6,6,6,6,6,6,6,6,0,0,0,0},
		'{6,6,6,6,6,6,6,6,0,0,0,0},
		'{6,6,6,6,6,6,6,6,0,0,0,0},
		'{6,6,6,6,6,6,6,6,0,0,0,0}};
		
		S_block_1 = '{
		'{6,6,6,6,0,0,0,0},
		'{6,6,6,6,0,0,0,0},
		'{6,6,6,6,0,0,0,0},
		'{6,6,6,6,0,0,0,0},
		'{6,6,6,6,6,6,6,6},
		'{6,6,6,6,6,6,6,6},
		'{6,6,6,6,6,6,6,6},
		'{6,6,6,6,6,6,6,6},
		'{0,0,0,0,6,6,6,6},
		'{0,0,0,0,6,6,6,6},
		'{0,0,0,0,6,6,6,6},
		'{0,0,0,0,6,6,6,6}};
		
		Z_block_0 = '{
		'{6,6,6,6,6,6,6,6,0,0,0,0},
		'{6,6,6,6,6,6,6,6,0,0,0,0},
		'{6,6,6,6,6,6,6,6,0,0,0,0},
		'{6,6,6,6,6,6,6,6,0,0,0,0},
		'{0,0,0,0,6,6,6,6,6,6,6,6},
		'{0,0,0,0,6,6,6,6,6,6,6,6},
		'{0,0,0,0,6,6,6,6,6,6,6,6},
		'{0,0,0,0,6,6,6,6,6,6,6,6}	};
		
		Z_block_1 = '{
		'{0,0,0,0,6,6,6,6},
		'{0,0,0,0,6,6,6,6},
		'{0,0,0,0,6,6,6,6},
		'{0,0,0,0,6,6,6,6},
		'{6,6,6,6,6,6,6,6},
		'{6,6,6,6,6,6,6,6},
		'{6,6,6,6,6,6,6,6},
		'{6,6,6,6,6,6,6,6},
		'{6,6,6,6,0,0,0,0},
		'{6,6,6,6,0,0,0,0},
		'{6,6,6,6,0,0,0,0},
		'{6,6,6,6,0,0,0,0}};
		
		T_block_0 = '{
		'{7,7,7,7,7,7,7,7,7,7,7,7},
		'{7,7,7,7,7,7,7,7,7,7,7,7},
		'{7,7,7,7,7,7,7,7,7,7,7,7},
		'{7,7,7,7,7,7,7,7,7,7,7,7},
		'{0,0,0,0,7,7,7,7,0,0,0,0},
		'{0,0,0,0,7,7,7,7,0,0,0,0},
		'{0,0,0,0,7,7,7,7,0,0,0,0},
		'{0,0,0,0,7,7,7,7,0,0,0,0}};
		
		T_block_1 = '{
		'{0,0,0,0,7,7,7,7},
		'{0,0,0,0,7,7,7,7},
		'{0,0,0,0,7,7,7,7},
		'{0,0,0,0,7,7,7,7},
		'{7,7,7,7,7,7,7,7},
		'{7,7,7,7,7,7,7,7},
		'{7,7,7,7,7,7,7,7},
		'{7,7,7,7,7,7,7,7},
		'{0,0,0,0,7,7,7,7},
		'{0,0,0,0,7,7,7,7},
		'{0,0,0,0,7,7,7,7},
		'{0,0,0,0,7,7,7,7}};
		
		T_block_2 = '{
		'{0,0,0,0,7,7,7,7,0,0,0,0},
		'{0,0,0,0,7,7,7,7,0,0,0,0},
		'{0,0,0,0,7,7,7,7,0,0,0,0},
		'{0,0,0,0,7,7,7,7,0,0,0,0},
		'{7,7,7,7,7,7,7,7,7,7,7,7},
		'{7,7,7,7,7,7,7,7,7,7,7,7},
		'{7,7,7,7,7,7,7,7,7,7,7,7},
		'{7,7,7,7,7,7,7,7,7,7,7,7}};
		
		T_block_3 = '{
		'{7,7,7,7,0,0,0,0},
		'{7,7,7,7,0,0,0,0},
		'{7,7,7,7,0,0,0,0},
		'{7,7,7,7,0,0,0,0},
		'{7,7,7,7,7,7,7,7},
		'{7,7,7,7,7,7,7,7},
		'{7,7,7,7,7,7,7,7},
		'{7,7,7,7,7,7,7,7},
		'{7,7,7,7,0,0,0,0},
		'{7,7,7,7,0,0,0,0},
		'{7,7,7,7,0,0,0,0},
		'{7,7,7,7,0,0,0,0}};

		TETRIS_h <= '{
		'{0,0,7,7,7,7,7,0,1,1,1,1,1,0,5,0,0,0,5,0,0,0,2,0,0,0,4,4,4,4,4,0,0,0,6,0,0,0,0,0},
		'{0,0,7,0,0,0,0,0,0,0,1,0,0,0,0,5,0,0,5,0,0,0,2,0,0,0,0,0,0,0,4,0,0,0,6,0,0,0,0,0},
		'{0,0,7,7,7,7,7,0,0,0,1,0,0,0,5,5,5,5,5,0,0,0,2,0,0,0,4,4,4,4,4,0,0,0,6,0,0,0,0,0},
		'{0,0,0,0,0,0,7,0,0,0,1,0,0,0,5,0,0,0,5,0,0,0,2,0,0,0,0,0,0,0,4,0,0,0,6,0,0,0,0,0},
		'{0,0,7,7,7,7,7,0,1,1,1,1,1,0,5,5,5,5,5,0,2,2,2,2,2,0,4,4,4,4,4,0,6,6,6,6,6,0,0,0}};
	
		game_over <= '{	
		'{0,4,0,0,0,4,0,6,6,6,6,6,0,0,0,8,0,0,0,1,1,1,1,1,0},
		'{0,0,4,0,0,4,0,0,0,0,0,6,0,8,8,0,8,8,0,1,0,0,0,1,0},
		'{0,4,4,4,4,4,0,6,6,6,6,6,0,8,0,0,0,8,0,1,0,0,0,1,0},
		'{0,4,0,0,0,4,0,0,0,0,0,6,0,8,0,0,0,8,0,1,0,0,0,1,0},
		'{0,4,4,4,4,4,0,6,6,6,6,6,0,8,0,0,0,8,0,1,1,1,1,1,0},
		'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
		'{0,5,5,5,5,5,0,2,0,0,0,2,0,4,0,0,0,4,0,6,6,6,6,6,0},
		'{0,0,0,0,0,5,0,2,0,0,0,2,0,4,0,0,0,4,0,6,0,0,0,6,0},
		'{0,5,5,5,5,5,0,2,0,2,0,2,0,4,4,4,4,4,0,6,6,0,0,6,0},
		'{0,0,0,0,0,5,0,2,2,0,2,2,0,4,0,0,0,4,0,0,0,0,0,6,0},
		'{0,5,5,5,5,5,0,2,0,0,0,2,0,4,4,4,4,4,0,6,6,6,6,6,0}};
		
		SCORE_Letters <= '{
		'{4,4,4,4,4,0,2,0,0,0,2,0,5,5,5,5,5,0,1,1,1,1,1,0,7,7,7,7,7},
		'{0,0,0,0,4,0,0,2,0,0,2,0,5,0,0,0,5,0,0,0,0,0,1,0,7,0,0,0,0},
		'{4,4,4,4,4,0,2,2,2,2,2,0,5,0,0,0,5,0,0,0,0,0,1,0,7,7,7,7,7},
		'{0,0,0,0,4,0,2,0,0,0,2,0,5,0,0,0,5,0,0,0,0,0,1,0,0,0,0,0,7},
		'{4,4,4,4,4,0,2,2,2,2,2,0,5,5,5,5,5,0,1,1,1,1,1,0,7,7,7,7,7}};
		
		zero <= '{
		'{9,9,9,9,9},
		'{9,0,0,0,9},
		'{9,0,0,0,9},
		'{9,0,0,0,9},
		'{9,9,9,9,9}};
		
		
		one <= '{
		'{0,0,9,0,0},
		'{0,0,9,0,0},
		'{0,0,9,0,0},
		'{0,0,9,0,0},
		'{0,0,9,0,0}};	
		
		two <= '{
		'{9,9,9,9,9},
		'{0,0,0,0,9},
		'{9,9,9,9,9},
		'{9,0,0,0,0},
		'{9,9,9,9,9}};

		three <= '{
		'{9,9,9,9,9},
		'{9,0,0,0,0},
		'{9,9,9,9,9},
		'{9,0,0,0,0},
		'{9,9,9,9,9}};
		
		
		
		four <= '{
		'{9,0,0,0,0},
		'{9,0,0,0,0},
		'{9,9,9,9,9},
		'{9,0,0,0,9},
		'{9,0,0,0,9}};
		
		five <= '{
		'{9,9,9,9,9},
		'{9,0,0,0,0},
		'{9,9,9,9,9},
		'{0,0,0,0,9},
		'{9,9,9,9,9}};
		
		six <= '{
		'{9,9,9,9,9},
		'{9,0,0,0,9},
		'{9,9,9,9,9},
		'{0,0,0,0,9},
		'{9,9,9,9,9}};
		
		seven <= '{
		'{9,0,0,0,0},
		'{9,0,0,0,0},
		'{9,0,0,0,0},
		'{9,0,0,0,9},
		'{9,9,9,9,9}};

		eight <= '{
		'{9,9,9,9,9},
		'{9,0,0,0,9},
		'{9,9,9,9,9},
		'{9,0,0,0,9},
		'{9,9,9,9,9}};	
		
		nine <= '{
		'{9,9,9,9,9},
		'{9,0,0,0,0},
		'{9,9,9,9,9},
		'{9,0,0,0,9},
		'{9,9,9,9,9}};
		
	 end
endmodule 